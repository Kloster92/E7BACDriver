** Profile: "Load step-Loadstep"  [ C:\Users\Jesper\Documents\GitHub\E7BACDriver\P-Spice\Simulering med 3f3\2. iteration\Flyback_2iteration_TEST-PSpiceFiles\Load step\Loadstep.sim ] 

** Creating circuit file "Loadstep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/Jesper/Documents/GitHub/E7BACDriver/P-Spice/Simulering med 3f3/uccx813-1.lib" 
.LIB "C:/Users/Jesper/Documents/GitHub/E7BACDriver/P-Spice/Simulering med 3f3/ntsv30120ctg.lib" 
.LIB "C:/Users/Jesper/Documents/GitHub/E7BACDriver/P-Spice/Simulering med 3f3/fdpf770n15a.lib" 
.LIB "C:/Cadence/SMPS PSpice Kursus/PSpice Files/Library/Smps/PSpice/Ferrite.lib" 
* From [PSPICE NETLIST] section of C:\Users\Jesper\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\pspice_demokit.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\sample_models.lib" 

*Analysis directives: 
.TRAN/OP 10ns 30ms 20ms 1us 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1.0u
.OPTIONS VNTOL= 10.0u
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Load step.net" 


.END
