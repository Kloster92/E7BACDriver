** Profile: "Gain-Phase-AC"  [ C:\Users\Nicolai Fransen\Documents\GitHub\E7BACDriver\P-Spice\Simulering med 3f3\Flyback_diagram TEST-PSpiceFiles\Gain-Phase\AC.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/Library/Smps/PSpice/Ferrite.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\pspice_demokit.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\sample_models.lib" 

*Analysis directives: 
.AC DEC 1000 10 100k
.STEP PARAM Pscale LIST 0.1 1 
.OPTIONS ADVCONV
.OPTIONS CONVAID
.OPTIONS METHOD= Default
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\Gain-Phase.net" 


.END
