** Profile: "Flyback_Linear-Tran"  [ C:\Users\Nicolai Fransen\Documents\GitHub\E7BACDriver\P-Spice\Simulering med 3f3\Flyback_E7BAC-PSpiceFiles\Flyback_Linear\Tran.sim ] 

** Creating circuit file "Tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../flyback_e7bac-pspicefiles/flyback_e7bac.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\pspice_demokit.lib" 
.lib "C:\Cadence\Company\OrCAD_PSpice\Models\sample_models.lib" 

*Analysis directives: 
.TRAN  0 1.1m 1m 10n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Flyback_Linear.net" 


.END
